--
-- File:   __PROJECT-NAME___tb.vhd
-- Author: __USER-NAME__
-- 
-- Created on __(format-time-string "%B %e, %Y, %l:%M %p")__
--

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity __PROJECT-NAME___tb is
end;

architecture __PROJECT-NAME___tb_arq of __PROJECT-NAME___tb is
begin
end;
