/**
 * File:   __PROJECT-NAME__.v
 * Author: __USER-NAME__
 * 
 * Created on __(format-time-string "%B %e, %Y, %l:%M %p")__
 */

module __PROJECT-NAME__ (/*PORTS*/);
endmodule // __PROJECT-NAME__
