--
-- File:   __PROJECT-NAME__.vhd
-- Author: __USER-NAME__
-- 
-- Created on __(format-time-string "%B %e, %Y, %l:%M %p")__
--

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity __PROJECT-NAME__ is
end;

architecture __PROJECT-NAME___arq of __PROJECT-NAME__ is
begin
end;
