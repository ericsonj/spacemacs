/**
 * File:   __PROJECT-NAME___tb.v
 * Author: __USER-NAME__
 * 
 * Created on __(format-time-string "%B %e, %Y, %l:%M %p")__
 */

module __PROJECT-NAME___tb (/**PORTS**/);
endmodule // __PROJECT-NAME___tb
